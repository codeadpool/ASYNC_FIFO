package afifo_tb_pkg;
  import uvm_pkg::*;
  
  `include "afifo_if.sv"
  `include "dut_harness.sv"
  `include "clkgen.sv"
endpackage
