package afifo_wr_agent_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "afifo_txn.sv"
  `include "afifo_wr_driver.svh"
  `include "afifo_wr_monitor.svh"
endpackage
